** Profile: "root-7"  [ E:\local\college\classes\2021bF\ECEN4013\ECEN4013\ADC\pspice\schematic\adc-pspicefiles\root\7.sim ] 

** Creating circuit file "7.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "E:\local\college\classes\2021bF\ECEN4013\ECEN4013\ADC\pspice\schematic\adc-pspicefiles\root\7\7_profile.inc" 
* Local Libraries :
.LIB "E:/local/college/classes/2021bF/ECEN4013/ECEN4013/ADC/pspice/models/cd4000.lib" 
.LIB "../../../adc-pspicefiles/adc.lib" 
.LIB "E:/local/college/classes/2021bF/ECEN4013/ECEN4013/ADC/pspice/models/tl082.lib" 
.LIB "E:/local/college/classes/2021bF/ECEN4013/ECEN4013/ADC/pspice/models/cd4066-cd4060/cd4066b.lib" 
.STMLIB "../../../adc-PSpiceFiles/ADC.stl" 
* From [PSPICE NETLIST] section of C:\Users\colli\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "E:\local\college\microg\saver2021\signals\pspice\models\Q50a02ch.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.3 0 
.OPTIONS ADVCONV
.OPTIONS DIGINITSTATE= 0
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\root.net" 


.END
