** Profile: "counter-counter"  [ E:\local\college\classes\2021bF\ECEN4013\ADC\circuits\schematic\adc-PSpiceFiles\counter\counter.sim ] 

** Creating circuit file "counter.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "E:\local\college\classes\2021bF\ECEN4013\ADC\circuits\schematic\adc-PSpiceFiles\counter\counter\counter_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\colli\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10u 0 10n 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\counter.net" 


.END
